///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: SE18_32
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbench();
`include "../Test/Test.v"
///////////////////////////////////////////////////////////////////////////////////
// Input: A (18-bit)
reg[17:0] A;
///////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
// Output: S (32-bit)
wire[31:0] S;
///////////////////////////////////////////////////////////////////////////////////

SE18_32 mySE(A, S);

initial begin
////////////////////////////////////////////////////////////////////////////////////////
// Test: Positive A
$display("Testing positive A=3782");
A=3782;   #10; 
////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////
// Test: Negative A
$display("Testing negative A=-43");
verifyEqual($signed(S), $signed(A));
////////////////////////////////////////////////////////////////////////////////////////

$display("All tests passed.");
end

endmodule
